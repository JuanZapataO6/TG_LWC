LIBRARY ieee;
USE ieee.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
USE ieee.numeric_std.ALL;
entity AesKey is
port (      
    En_In   : in std_logic; -- Flag for start FMS
    Ena_Out : out std_logic;
    Clk : in std_logic; -- Clock signal 
    --Read Memory bank of key from DataGenerate 
    Rd_En_K : out std_logic;
    Data_in_K : in std_logic_vector (7 downto 0);  
    Addr_Rd_K : out std_logic_vector (3 DOWNTO 0);
    --Output Memory Bank yourself
    Rd_En_eK : in std_logic;
    Addr_Rd_eK : in std_logic_vector (5 DOWNTO 0);
    Data_Out_eK : out std_logic_vector (31 downto 0) 
);
end AesKey;
architecture RTL of AesKey is
component MemBnk
    generic(    
        w:integer;--width of word
        d:integer;--Numbers of words 
        a:integer --width of Address
    );
    port( 
        Wr_En    : in  std_logic;
        Rd_En    : in  std_logic;        
        Rst      : in  std_logic;
        Clk      : in  std_logic;
        Addr_In  : in  std_logic_vector (a-1 downto 0);
        Addr_Out : in  std_logic_vector (a-1 downto 0);
        Data_in  : in  std_logic_vector (w-1 downto 0);
        Data_Out : out std_logic_vector (w-1 downto 0)
    );
end component; 
component Register_A
    generic(
        w:integer--width of word
    );
    port (
        DD_IN  : in  std_logic_vector (w-1 downto 0);
        DD_OUT : out std_logic_vector (w-1 downto 0);
        Clk    : in  std_logic
    );
end component Register_A;
TYPE estado is (s0, s1,s2,s3,s4,s5,s6,s7,s8,s9,s10,s11,s12,s13,s14,s15,s16,s17,s18,s19,s20);
SIGNAL presente:estado:=s0;
--signals for write in memory bank hear
signal Wr_En_eK : std_logic;
signal Rst  : std_logic;
signal Addr_Wr_eK : std_logic_vector (5 downto 0);
signal Data_In_eK : std_logic_vector (31 downto 0);
signal Data_Rin_K : std_logic_vector (7 downto 0);  
begin 
--Component for AesKey Places for 32 bits 
uRin_K :  Register_A 
    generic map (
        w => 8
    ) 
    Port map (
    DD_IN  => Data_In_K,
    DD_OUT => Data_RIn_K,
    Clk    => clk
    );
uEkey: MemBnk
    generic map(
        w => 32, --Witdth of words
        d => 44, --Numbers of Words
        a => 6   --Witdth of Address
    )
    Port Map (  
        Wr_En    => Wr_En_eK,   --signal 
        Rd_En    => Rd_En_eK,   --port 
        Rst      => Rst,        --signal 
        Clk      => clk,        --port
        Addr_In  => Addr_Wr_eK, --signal 
        Addr_Out => Addr_Rd_eK, --port
        Data_in  => Data_In_eK, --signal 
        Data_Out => Data_Out_eK --port
    );
STat: process (clk,presente)
type word is array (0 to 43) of std_logic_vector (31 downto 0);
variable eKeyAux : word;
type C_M0 is array (0 to 255) of std_logic_vector (31 downto 0);
constant M0 : C_M0:= (
    x"a56363c6", x"847c7cf8", x"997777ee", x"8d7b7bf6", x"0df2f2ff", x"bd6b6bd6", x"b16f6fde", x"54c5c591",
    x"50303060", x"03010102", x"a96767ce", x"7d2b2b56", x"19fefee7", x"62d7d7b5", x"e6abab4d", x"9a7676ec",
    x"45caca8f", x"9d82821f", x"40c9c989", x"877d7dfa", x"15fafaef", x"eb5959b2", x"c947478e", x"0bf0f0fb",
    x"ecadad41", x"67d4d4b3", x"fda2a25f", x"eaafaf45", x"bf9c9c23", x"f7a4a453", x"967272e4", x"5bc0c09b",
    x"c2b7b775", x"1cfdfde1", x"ae93933d", x"6a26264c", x"5a36366c", x"413f3f7e", x"02f7f7f5", x"4fcccc83",
    x"5c343468", x"f4a5a551", x"34e5e5d1", x"08f1f1f9", x"937171e2", x"73d8d8ab", x"53313162", x"3f15152a",
    x"0c040408", x"52c7c795", x"65232346", x"5ec3c39d", x"28181830", x"a1969637", x"0f05050a", x"b59a9a2f",
    x"0907070e", x"36121224", x"9b80801b", x"3de2e2df", x"26ebebcd", x"6927274e", x"cdb2b27f", x"9f7575ea",
    x"1b090912", x"9e83831d", x"742c2c58", x"2e1a1a34", x"2d1b1b36", x"b26e6edc", x"ee5a5ab4", x"fba0a05b",
    x"f65252a4", x"4d3b3b76", x"61d6d6b7", x"ceb3b37d", x"7b292952", x"3ee3e3dd", x"712f2f5e", x"97848413",
    x"f55353a6", x"68d1d1b9", x"00000000", x"2cededc1", x"60202040", x"1ffcfce3", x"c8b1b179", x"ed5b5bb6",
    x"be6a6ad4", x"46cbcb8d", x"d9bebe67", x"4b393972", x"de4a4a94", x"d44c4c98", x"e85858b0", x"4acfcf85",
    x"6bd0d0bb", x"2aefefc5", x"e5aaaa4f", x"16fbfbed", x"c5434386", x"d74d4d9a", x"55333366", x"94858511",
    x"cf45458a", x"10f9f9e9", x"06020204", x"817f7ffe", x"f05050a0", x"443c3c78", x"ba9f9f25", x"e3a8a84b",
    x"f35151a2", x"fea3a35d", x"c0404080", x"8a8f8f05", x"ad92923f", x"bc9d9d21", x"48383870", x"04f5f5f1",
    x"dfbcbc63", x"c1b6b677", x"75dadaaf", x"63212142", x"30101020", x"1affffe5", x"0ef3f3fd", x"6dd2d2bf",
    x"4ccdcd81", x"140c0c18", x"35131326", x"2fececc3", x"e15f5fbe", x"a2979735", x"cc444488", x"3917172e",
    x"57c4c493", x"f2a7a755", x"827e7efc", x"473d3d7a", x"ac6464c8", x"e75d5dba", x"2b191932", x"957373e6",
    x"a06060c0", x"98818119", x"d14f4f9e", x"7fdcdca3", x"66222244", x"7e2a2a54", x"ab90903b", x"8388880b",
    x"ca46468c", x"29eeeec7", x"d3b8b86b", x"3c141428", x"79dedea7", x"e25e5ebc", x"1d0b0b16", x"76dbdbad",
    x"3be0e0db", x"56323264", x"4e3a3a74", x"1e0a0a14", x"db494992", x"0a06060c", x"6c242448", x"e45c5cb8",
    x"5dc2c29f", x"6ed3d3bd", x"efacac43", x"a66262c4", x"a8919139", x"a4959531", x"37e4e4d3", x"8b7979f2",
    x"32e7e7d5", x"43c8c88b", x"5937376e", x"b76d6dda", x"8c8d8d01", x"64d5d5b1", x"d24e4e9c", x"e0a9a949",
    x"b46c6cd8", x"fa5656ac", x"07f4f4f3", x"25eaeacf", x"af6565ca", x"8e7a7af4", x"e9aeae47", x"18080810",
    x"d5baba6f", x"887878f0", x"6f25254a", x"722e2e5c", x"241c1c38", x"f1a6a657", x"c7b4b473", x"51c6c697",
    x"23e8e8cb", x"7cdddda1", x"9c7474e8", x"211f1f3e", x"dd4b4b96", x"dcbdbd61", x"868b8b0d", x"858a8a0f",
    x"907070e0", x"423e3e7c", x"c4b5b571", x"aa6666cc", x"d8484890", x"05030306", x"01f6f6f7", x"120e0e1c",
    x"a36161c2", x"5f35356a", x"f95757ae", x"d0b9b969", x"91868617", x"58c1c199", x"271d1d3a", x"b99e9e27",
    x"38e1e1d9", x"13f8f8eb", x"b398982b", x"33111122", x"bb6969d2", x"70d9d9a9", x"898e8e07", x"a7949433",
    x"b69b9b2d", x"221e1e3c", x"92878715", x"20e9e9c9", x"49cece87", x"ff5555aa", x"78282850", x"7adfdfa5",
    x"8f8c8c03", x"f8a1a159", x"80898909", x"170d0d1a", x"dabfbf65", x"31e6e6d7", x"c6424284", x"b86868d0",
    x"c3414182", x"b0999929", x"772d2d5a", x"110f0f1e", x"cbb0b07b", x"fc5454a8", x"d6bbbb6d", x"3a16162c"
);
type C_M1 is array (0 to 255) of std_logic_vector (31 downto 0);
constant M1 : C_M1:= (
    x"6363c6a5", x"7c7cf884", x"7777ee99", x"7b7bf68d", x"f2f2ff0d", x"6b6bd6bd", x"6f6fdeb1", x"c5c59154", 
    x"30306050", x"01010203", x"6767cea9", x"2b2b567d", x"fefee719", x"d7d7b562", x"abab4de6", x"7676ec9a", 
    x"caca8f45", x"82821f9d", x"c9c98940", x"7d7dfa87", x"fafaef15", x"5959b2eb", x"47478ec9", x"f0f0fb0b", 
    x"adad41ec", x"d4d4b367", x"a2a25ffd", x"afaf45ea", x"9c9c23bf", x"a4a453f7", x"7272e496", x"c0c09b5b", 
    x"b7b775c2", x"fdfde11c", x"93933dae", x"26264c6a", x"36366c5a", x"3f3f7e41", x"f7f7f502", x"cccc834f", 
    x"3434685c", x"a5a551f4", x"e5e5d134", x"f1f1f908", x"7171e293", x"d8d8ab73", x"31316253", x"15152a3f", 
    x"0404080c", x"c7c79552", x"23234665", x"c3c39d5e", x"18183028", x"969637a1", x"05050a0f", x"9a9a2fb5", 
    x"07070e09", x"12122436", x"80801b9b", x"e2e2df3d", x"ebebcd26", x"27274e69", x"b2b27fcd", x"7575ea9f", 
    x"0909121b", x"83831d9e", x"2c2c5874", x"1a1a342e", x"1b1b362d", x"6e6edcb2", x"5a5ab4ee", x"a0a05bfb", 
    x"5252a4f6", x"3b3b764d", x"d6d6b761", x"b3b37dce", x"2929527b", x"e3e3dd3e", x"2f2f5e71", x"84841397", 
    x"5353a6f5", x"d1d1b968", x"00000000", x"ededc12c", x"20204060", x"fcfce31f", x"b1b179c8", x"5b5bb6ed", 
    x"6a6ad4be", x"cbcb8d46", x"bebe67d9", x"3939724b", x"4a4a94de", x"4c4c98d4", x"5858b0e8", x"cfcf854a", 
    x"d0d0bb6b", x"efefc52a", x"aaaa4fe5", x"fbfbed16", x"434386c5", x"4d4d9ad7", x"33336655", x"85851194", 
    x"45458acf", x"f9f9e910", x"02020406", x"7f7ffe81", x"5050a0f0", x"3c3c7844", x"9f9f25ba", x"a8a84be3", 
    x"5151a2f3", x"a3a35dfe", x"404080c0", x"8f8f058a", x"92923fad", x"9d9d21bc", x"38387048", x"f5f5f104", 
    x"bcbc63df", x"b6b677c1", x"dadaaf75", x"21214263", x"10102030", x"ffffe51a", x"f3f3fd0e", x"d2d2bf6d", 
    x"cdcd814c", x"0c0c1814", x"13132635", x"ececc32f", x"5f5fbee1", x"979735a2", x"444488cc", x"17172e39", 
    x"c4c49357", x"a7a755f2", x"7e7efc82", x"3d3d7a47", x"6464c8ac", x"5d5dbae7", x"1919322b", x"7373e695", 
    x"6060c0a0", x"81811998", x"4f4f9ed1", x"dcdca37f", x"22224466", x"2a2a547e", x"90903bab", x"88880b83", 
    x"46468cca", x"eeeec729", x"b8b86bd3", x"1414283c", x"dedea779", x"5e5ebce2", x"0b0b161d", x"dbdbad76", 
    x"e0e0db3b", x"32326456", x"3a3a744e", x"0a0a141e", x"494992db", x"06060c0a", x"2424486c", x"5c5cb8e4", 
    x"c2c29f5d", x"d3d3bd6e", x"acac43ef", x"6262c4a6", x"919139a8", x"959531a4", x"e4e4d337", x"7979f28b", 
    x"e7e7d532", x"c8c88b43", x"37376e59", x"6d6ddab7", x"8d8d018c", x"d5d5b164", x"4e4e9cd2", x"a9a949e0", 
    x"6c6cd8b4", x"5656acfa", x"f4f4f307", x"eaeacf25", x"6565caaf", x"7a7af48e", x"aeae47e9", x"08081018", 
    x"baba6fd5", x"7878f088", x"25254a6f", x"2e2e5c72", x"1c1c3824", x"a6a657f1", x"b4b473c7", x"c6c69751", 
    x"e8e8cb23", x"dddda17c", x"7474e89c", x"1f1f3e21", x"4b4b96dd", x"bdbd61dc", x"8b8b0d86", x"8a8a0f85", 
    x"7070e090", x"3e3e7c42", x"b5b571c4", x"6666ccaa", x"484890d8", x"03030605", x"f6f6f701", x"0e0e1c12", 
    x"6161c2a3", x"35356a5f", x"5757aef9", x"b9b969d0", x"86861791", x"c1c19958", x"1d1d3a27", x"9e9e27b9", 
    x"e1e1d938", x"f8f8eb13", x"98982bb3", x"11112233", x"6969d2bb", x"d9d9a970", x"8e8e0789", x"949433a7", 
    x"9b9b2db6", x"1e1e3c22", x"87871592", x"e9e9c920", x"cece8749", x"5555aaff", x"28285078", x"dfdfa57a", 
    x"8c8c038f", x"a1a159f8", x"89890980", x"0d0d1a17", x"bfbf65da", x"e6e6d731", x"424284c6", x"6868d0b8", 
    x"414182c3", x"999929b0", x"2d2d5a77", x"0f0f1e11", x"b0b07bcb", x"5454a8fc", x"bbbb6dd6", x"16162c3a"
);
type C_M2 is array (0 to 255) of std_logic_vector (31 downto 0);
constant M2 : C_M2:= (
    x"63c6a563", x"7cf8847c", x"77ee9977", x"7bf68d7b", x"f2ff0df2", x"6bd6bd6b", x"6fdeb16f", x"c59154c5", 
    x"30605030", x"01020301", x"67cea967", x"2b567d2b", x"fee719fe", x"d7b562d7", x"ab4de6ab", x"76ec9a76", 
    x"ca8f45ca", x"821f9d82", x"c98940c9", x"7dfa877d", x"faef15fa", x"59b2eb59", x"478ec947", x"f0fb0bf0", 
    x"ad41ecad", x"d4b367d4", x"a25ffda2", x"af45eaaf", x"9c23bf9c", x"a453f7a4", x"72e49672", x"c09b5bc0", 
    x"b775c2b7", x"fde11cfd", x"933dae93", x"264c6a26", x"366c5a36", x"3f7e413f", x"f7f502f7", x"cc834fcc", 
    x"34685c34", x"a551f4a5", x"e5d134e5", x"f1f908f1", x"71e29371", x"d8ab73d8", x"31625331", x"152a3f15", 
    x"04080c04", x"c79552c7", x"23466523", x"c39d5ec3", x"18302818", x"9637a196", x"050a0f05", x"9a2fb59a", 
    x"070e0907", x"12243612", x"801b9b80", x"e2df3de2", x"ebcd26eb", x"274e6927", x"b27fcdb2", x"75ea9f75", 
    x"09121b09", x"831d9e83", x"2c58742c", x"1a342e1a", x"1b362d1b", x"6edcb26e", x"5ab4ee5a", x"a05bfba0", 
    x"52a4f652", x"3b764d3b", x"d6b761d6", x"b37dceb3", x"29527b29", x"e3dd3ee3", x"2f5e712f", x"84139784", 
    x"53a6f553", x"d1b968d1", x"00000000", x"edc12ced", x"20406020", x"fce31ffc", x"b179c8b1", x"5bb6ed5b", 
    x"6ad4be6a", x"cb8d46cb", x"be67d9be", x"39724b39", x"4a94de4a", x"4c98d44c", x"58b0e858", x"cf854acf", 
    x"d0bb6bd0", x"efc52aef", x"aa4fe5aa", x"fbed16fb", x"4386c543", x"4d9ad74d", x"33665533", x"85119485", 
    x"458acf45", x"f9e910f9", x"02040602", x"7ffe817f", x"50a0f050", x"3c78443c", x"9f25ba9f", x"a84be3a8", 
    x"51a2f351", x"a35dfea3", x"4080c040", x"8f058a8f", x"923fad92", x"9d21bc9d", x"38704838", x"f5f104f5", 
    x"bc63dfbc", x"b677c1b6", x"daaf75da", x"21426321", x"10203010", x"ffe51aff", x"f3fd0ef3", x"d2bf6dd2", 
    x"cd814ccd", x"0c18140c", x"13263513", x"ecc32fec", x"5fbee15f", x"9735a297", x"4488cc44", x"172e3917", 
    x"c49357c4", x"a755f2a7", x"7efc827e", x"3d7a473d", x"64c8ac64", x"5dbae75d", x"19322b19", x"73e69573", 
    x"60c0a060", x"81199881", x"4f9ed14f", x"dca37fdc", x"22446622", x"2a547e2a", x"903bab90", x"880b8388", 
    x"468cca46", x"eec729ee", x"b86bd3b8", x"14283c14", x"dea779de", x"5ebce25e", x"0b161d0b", x"dbad76db", 
    x"e0db3be0", x"32645632", x"3a744e3a", x"0a141e0a", x"4992db49", x"060c0a06", x"24486c24", x"5cb8e45c", 
    x"c29f5dc2", x"d3bd6ed3", x"ac43efac", x"62c4a662", x"9139a891", x"9531a495", x"e4d337e4", x"79f28b79", 
    x"e7d532e7", x"c88b43c8", x"376e5937", x"6ddab76d", x"8d018c8d", x"d5b164d5", x"4e9cd24e", x"a949e0a9", 
    x"6cd8b46c", x"56acfa56", x"f4f307f4", x"eacf25ea", x"65caaf65", x"7af48e7a", x"ae47e9ae", x"08101808", 
    x"ba6fd5ba", x"78f08878", x"254a6f25", x"2e5c722e", x"1c38241c", x"a657f1a6", x"b473c7b4", x"c69751c6", 
    x"e8cb23e8", x"dda17cdd", x"74e89c74", x"1f3e211f", x"4b96dd4b", x"bd61dcbd", x"8b0d868b", x"8a0f858a", 
    x"70e09070", x"3e7c423e", x"b571c4b5", x"66ccaa66", x"4890d848", x"03060503", x"f6f701f6", x"0e1c120e", 
    x"61c2a361", x"356a5f35", x"57aef957", x"b969d0b9", x"86179186", x"c19958c1", x"1d3a271d", x"9e27b99e", 
    x"e1d938e1", x"f8eb13f8", x"982bb398", x"11223311", x"69d2bb69", x"d9a970d9", x"8e07898e", x"9433a794", 
    x"9b2db69b", x"1e3c221e", x"87159287", x"e9c920e9", x"ce8749ce", x"55aaff55", x"28507828", x"dfa57adf", 
    x"8c038f8c", x"a159f8a1", x"89098089", x"0d1a170d", x"bf65dabf", x"e6d731e6", x"4284c642", x"68d0b868", 
    x"4182c341", x"9929b099", x"2d5a772d", x"0f1e110f", x"b07bcbb0", x"54a8fc54", x"bb6dd6bb", x"162c3a16"
);
type C_M3 is array (0 to 255) of std_logic_vector (31 downto 0);
constant M3 : C_M3:= (
    x"c6a56363", x"f8847c7c", x"ee997777", x"f68d7b7b", x"ff0df2f2", x"d6bd6b6b", x"deb16f6f", x"9154c5c5", 
    x"60503030", x"02030101", x"cea96767", x"567d2b2b", x"e719fefe", x"b562d7d7", x"4de6abab", x"ec9a7676", 
    x"8f45caca", x"1f9d8282", x"8940c9c9", x"fa877d7d", x"ef15fafa", x"b2eb5959", x"8ec94747", x"fb0bf0f0", 
    x"41ecadad", x"b367d4d4", x"5ffda2a2", x"45eaafaf", x"23bf9c9c", x"53f7a4a4", x"e4967272", x"9b5bc0c0", 
    x"75c2b7b7", x"e11cfdfd", x"3dae9393", x"4c6a2626", x"6c5a3636", x"7e413f3f", x"f502f7f7", x"834fcccc", 
    x"685c3434", x"51f4a5a5", x"d134e5e5", x"f908f1f1", x"e2937171", x"ab73d8d8", x"62533131", x"2a3f1515", 
    x"080c0404", x"9552c7c7", x"46652323", x"9d5ec3c3", x"30281818", x"37a19696", x"0a0f0505", x"2fb59a9a", 
    x"0e090707", x"24361212", x"1b9b8080", x"df3de2e2", x"cd26ebeb", x"4e692727", x"7fcdb2b2", x"ea9f7575", 
    x"121b0909", x"1d9e8383", x"58742c2c", x"342e1a1a", x"362d1b1b", x"dcb26e6e", x"b4ee5a5a", x"5bfba0a0", 
    x"a4f65252", x"764d3b3b", x"b761d6d6", x"7dceb3b3", x"527b2929", x"dd3ee3e3", x"5e712f2f", x"13978484", 
    x"a6f55353", x"b968d1d1", x"00000000", x"c12ceded", x"40602020", x"e31ffcfc", x"79c8b1b1", x"b6ed5b5b", 
    x"d4be6a6a", x"8d46cbcb", x"67d9bebe", x"724b3939", x"94de4a4a", x"98d44c4c", x"b0e85858", x"854acfcf", 
    x"bb6bd0d0", x"c52aefef", x"4fe5aaaa", x"ed16fbfb", x"86c54343", x"9ad74d4d", x"66553333", x"11948585", 
    x"8acf4545", x"e910f9f9", x"04060202", x"fe817f7f", x"a0f05050", x"78443c3c", x"25ba9f9f", x"4be3a8a8", 
    x"a2f35151", x"5dfea3a3", x"80c04040", x"058a8f8f", x"3fad9292", x"21bc9d9d", x"70483838", x"f104f5f5", 
    x"63dfbcbc", x"77c1b6b6", x"af75dada", x"42632121", x"20301010", x"e51affff", x"fd0ef3f3", x"bf6dd2d2", 
    x"814ccdcd", x"18140c0c", x"26351313", x"c32fecec", x"bee15f5f", x"35a29797", x"88cc4444", x"2e391717", 
    x"9357c4c4", x"55f2a7a7", x"fc827e7e", x"7a473d3d", x"c8ac6464", x"bae75d5d", x"322b1919", x"e6957373", 
    x"c0a06060", x"19988181", x"9ed14f4f", x"a37fdcdc", x"44662222", x"547e2a2a", x"3bab9090", x"0b838888", 
    x"8cca4646", x"c729eeee", x"6bd3b8b8", x"283c1414", x"a779dede", x"bce25e5e", x"161d0b0b", x"ad76dbdb", 
    x"db3be0e0", x"64563232", x"744e3a3a", x"141e0a0a", x"92db4949", x"0c0a0606", x"486c2424", x"b8e45c5c", 
    x"9f5dc2c2", x"bd6ed3d3", x"43efacac", x"c4a66262", x"39a89191", x"31a49595", x"d337e4e4", x"f28b7979", 
    x"d532e7e7", x"8b43c8c8", x"6e593737", x"dab76d6d", x"018c8d8d", x"b164d5d5", x"9cd24e4e", x"49e0a9a9", 
    x"d8b46c6c", x"acfa5656", x"f307f4f4", x"cf25eaea", x"caaf6565", x"f48e7a7a", x"47e9aeae", x"10180808", 
    x"6fd5baba", x"f0887878", x"4a6f2525", x"5c722e2e", x"38241c1c", x"57f1a6a6", x"73c7b4b4", x"9751c6c6", 
    x"cb23e8e8", x"a17cdddd", x"e89c7474", x"3e211f1f", x"96dd4b4b", x"61dcbdbd", x"0d868b8b", x"0f858a8a", 
    x"e0907070", x"7c423e3e", x"71c4b5b5", x"ccaa6666", x"90d84848", x"06050303", x"f701f6f6", x"1c120e0e", 
    x"c2a36161", x"6a5f3535", x"aef95757", x"69d0b9b9", x"17918686", x"9958c1c1", x"3a271d1d", x"27b99e9e", 
    x"d938e1e1", x"eb13f8f8", x"2bb39898", x"22331111", x"d2bb6969", x"a970d9d9", x"07898e8e", x"33a79494", 
    x"2db69b9b", x"3c221e1e", x"15928787", x"c920e9e9", x"8749cece", x"aaff5555", x"50782828", x"a57adfdf", 
    x"038f8c8c", x"59f8a1a1", x"09808989", x"1a170d0d", x"65dabfbf", x"d731e6e6", x"84c64242", x"d0b86868", 
    x"82c34141", x"29b09999", x"5a772d2d", x"1e110f0f", x"7bcbb0b0", x"a8fc5454", x"6dd6bbbb", x"2c3a1616"
);
variable Finish_En  : std_logic:= '0';
variable Finish_No  : std_logic:= '0';
variable Addr_Aux   : std_logic_vector (5 downto 0) := "000000";      
variable Addr_Aux_eK   : std_logic_vector (5 downto 0) := "000000";
begin 
if clk 'event and clk = '1' then
    if En_In = '1' then 
        case presente is
            when s0 =>
                presente <= s1;
                Rd_En_K <= '0';
                --Addr_Aux := Addr_Aux + 1; 
                Addr_Rd_K <= Addr_Aux(Addr_Aux'length-3 downto 0);
                Data_In_eK <= M0(to_integer(unsigned(Addr_Aux)));
            when s1 => 
                presente <= s2;
                Rd_En_K <= '0';
                Addr_Aux := Addr_Aux + 1; 
                Addr_Rd_K <= Addr_Aux(Addr_Aux'length-3 downto 0);
                Data_In_eK <= M0(to_integer(unsigned(Addr_Aux)));
                --Data_In_eK <= x"000000" & Data_Rin_K;
            when s2 => 
                presente <= s3;
                Rd_En_K <= '0';
                Addr_Aux := Addr_Aux + 1; 
                Addr_Rd_K <= Addr_Aux(Addr_Aux'length-3 downto 0);
                Data_In_eK <= M0(to_integer(unsigned(Addr_Aux)));
            when s3 => 
                presente <= s4;
                Rd_En_K <= '0';
                Addr_Aux := Addr_Aux + 1; 
                Addr_Rd_K <= Addr_Aux(Addr_Aux'length-3 downto 0);
                Data_In_eK <= x"000000" & Data_Rin_K;
                
            when s4 => 
                presente <= s5;
                Rd_En_K <= '0';
                --Addr_Aux := Addr_Aux + 1; 
                Addr_Rd_K <= Addr_Aux(Addr_Aux'length-3 downto 0);
                Data_In_eK <= x"0000" & Data_Rin_K & Data_In_eK(7 downto 0);
            when s5 => 
                presente <= s6;
                Rd_En_K <= '0';
                --Addr_Aux := Addr_Aux + 1; 
                Addr_Rd_K <= Addr_Aux(Addr_Aux'length-3 downto 0);
                Data_In_eK <= x"00" & Data_Rin_K & Data_In_eK(15 downto 0);
            when s6 => 
                presente <= s7;
                Rd_En_K <= '1';
                --Addr_Aux := Addr_Aux + 1; 
                Addr_Rd_K <= Addr_Aux(Addr_Aux'length-3 downto 0);
                Data_In_eK <= Data_Rin_K & Data_In_eK(23 downto 0);
            when s7 => 
                presente <= s8;
                Rd_En_K <= '1';
                Wr_En_eK <= '0';
                eKeyAux(to_integer(unsigned(Addr_Aux_eK))) := Data_In_eK; 
                Addr_Wr_eK <= Addr_Aux_eK;
                Addr_Aux := Addr_Aux + 1; 
                Addr_Rd_K <= Addr_Aux(Addr_Aux'length-3 downto 0);
            when s8 => 
                if Addr_Aux_eK = "000011" then  
                    presente <= s9;
                else
                    presente <= s0;
                end if;
                Rd_En_K <= '1';
                Wr_En_eK <= '1';
                Addr_Aux_eK := Addr_Aux_eK + 1; 
                Addr_Rd_K <= Addr_Aux(Addr_Aux'length-3 downto 0);
            when s9 => 
                presente <= s10;
                Data_In_eK <= eKeyAux(to_integer(unsigned(Addr_Aux_eK - 4))) ;
            when others => null;
        end case;
    end if;
end if;
end process;
end RTL;